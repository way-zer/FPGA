module Root (
    input clkI,
    output [7:0] rowO,colR,colG//点阵输出接口
);
    Matrix m1(clkI,{
        2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b10,
        2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,
        2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,
        2'b00,2'b00,2'b00,2'b00,2'b11,2'b00,2'b00,2'b00,
        2'b00,2'b00,2'b00,2'b11,2'b00,2'b00,2'b00,2'b00,
        2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,
        2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,
        2'b01,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00,2'b00
    },rowO,colR,colG);
endmodule